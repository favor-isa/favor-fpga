`default_nettype none

module top_sim(
    input wire i_clk
);

endmodule