/* verilator lint_off UNUSEDSIGNAL */
module decoder(
    input wire        i_clk,
    input wire [31:0] i_insn,
    output reg        o_valid = 0,
    output reg        o_halt = 0
);

// The "kind" of instruction.
wire [1:0] k;

// K0 instruction identifier.
wire [3:0] k0;

// Singleton instruction identifier.
wire [24:0] sng;

assign k   = i_insn[30:29];
assign k0  = i_insn[28:25];
assign sng = i_insn[24:0];

`include "cpustate.vinc"

// Handle singleton instructions.
always @(posedge i_clk) if(k == 2'b00 && k0 == 4'b0000) begin
    o_valid <= 1;
    case(sng)
        25'b0: o_halt <= 1;
        default: o_valid <= 0;
    endcase
end

always @(posedge i_clk) if(k != 2'b00) begin
    o_valid <= 0;
end

// always @(posedge i_clk) begin
//     o_valid <= 0;

//     case(k)
//         2'b00: begin
//             case(k0)
//                 2'b00: begin

//                 end

//             endcase
//         end
//         2'b01: begin
//         end
//         2'b10: begin
//         end
//         2'b11: begin
//         end
//     endcase
// end

endmodule
